// Code your design here
module AND_gate(input wire a, input wire b, output wire out);
  
  assign out = (a & b);
  
endmodule