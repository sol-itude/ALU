// Code your design here
module AND_gate(input a,b, output out);
  
  assign out = (a & b);
  
endmodule